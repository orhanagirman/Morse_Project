module adcproject2(output a,b,c,d,e,f,g,q0,w0,e0,q1,w1,e1,q2,w2,e2, input i7,i6,i5,i4,i3,i2,ia,i0);

wire p0,g0,f0,p1,g1,f1,p2,g2,f2;

binarycomparator aa(p0,g0,f0,0,1,0,i3,i2,ia,i0,0,1,1,1);
binarycomparator ab(q0,w0,e0,p0,g0,f0,i7,i6,i5,i4,0,0,1,0);

binarycomparator ac(p1,g1,f1,0,1,0,i3,i2,ia,i0,0,1,0,0);
binarycomparator ad(q1,w1,e1,p1,g1,f1,i7,i6,i5,i4,0,1,1,1);

binarycomparator ae(p2,g2,f2,0,1,0,i3,i2,ia,i0,0,0,1,0);
binarycomparator af(q2,w2,e2,p2,g2,f2,i7,i6,i5,i4,1,1,0,0);

assign a = ~((q0&~w0&~e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&~w2&e2));
assign b = ~((q0&~w0&~e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&w0&~e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&~w2&e2));
assign c = ~((q0&~w0&~e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&w0&~e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&~w2&e2));
assign d = ~((q0&~w0&~e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&~w2&e2));
assign e = ~((q0&~w0&~e0&q1&~w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&q2&~w2&~e2));
assign f = ~(q0&~w0&~e0&q1&~w1&~e1&q2&~w2&~e2);
assign g = ~((~q0&~w0&e0&~q1&w1&~e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&q2&~w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&w2&~e2)|(~q0&~w0&e0&~q1&~w1&e1&~q2&~w2&e2));

endmodule



module binarycomparator (output K,L,M, input x,y,z,A3,A2,A1,A0,B3,B2,B1,B0);


assign K = (x&~y&~z&~A3&B3)|(~x&y&~z&~A3&B3)|(~x&~y&z&~A3&B3)|((x&~y&~z)&((A3|~B3)&(~A3|B3))&(~A2&B2))|((~x&y&~z)&((A3|~B3)&(~A3|B3))&(~A2&B2))|((~x&~y&z)&((A3|~B3)&(~A3|B3))&(~A2&B2))|((x&~y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&(~A1&B1))|((~x&y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&(~A1&B1))|((~x&~y&z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&(~A1&B1))|((x&~y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&(~A0&B0))|((~x&y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&(~A0&B0))|((~x&~y&z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&(~A0&B0))|((x&~y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&((A0|~B0)&(~A0|B0)));
assign L = ((~x&y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&((A0|~B0)&(~A0|B0)));
assign M = (x&~y&~z&A3&~B3)|(~x&y&~z&A3&~B3)|(~x&~y&z&A3&~B3)|((x&~y&~z)&((A3|~B3)&(~A3|B3))&(A2&~B2))|((~x&y&~z)&((A3|~B3)&(~A3|B3))&(A2&~B2))|((~x&~y&z)&((A3|~B3)&(~A3|B3))&(A2&~B2))|((x&~y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&(A1&~B1))|((~x&y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&(A1&~B1))|((~x&~y&z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&(A1&~B1))|((x&~y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&(A0&~B0))|((~x&y&~z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&(A0&~B0))|((~x&~y&z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&(A0&~B0))|((~x&~y&z)&((A3|~B3)&(~A3|B3))&((A2|~B2)&(~A2|B2))&((A1|~B1)&(~A1|B1))&((A0|~B0)&(~A0|B0)));

endmodule
